 
module AND_gate (a, b, c);
  input a, b;
  output c;
  wire a, b, c;
  assign c = a & b;
endmodule