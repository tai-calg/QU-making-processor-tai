module inst_decoder(
    input [1:0] alu_op,
    input [2:0] funct3,
    input funct7b5,
    output wire [3:0] alu_ctrl,
    output wire [1:0] byte_size,
    output wire [1:0] sgn_ext_src,
    output wire rd2ext_src
);


    function [8:0] inst_decode_fn(
        input [1:0] alu_op,
        input [2:0] funct3,
        input funct7b5
    );
        /// output = 9'b aluctrl_bytesize_sgnextsrc_rd2extsrc
        begin
            case (alu_op)
                2'b00: begin // Load
                    case (funct3) 
                        3'b000: inst_decode_fn = 9'b0000_10_01_0; //1byte load(lb)
                        3'b001: inst_decode_fn = 9'b0000_01_10_0; //2byte load(lh)
                        3'b010: inst_decode_fn = 9'b0000_00_00_0; //4byte load(lw)
                        3'b100: inst_decode_fn = 9'b0000_10_00_0; //1byte load(lbu)
                    endcase
                end
                2'b01: begin // Branch
                    case (funct3) 
                        3'b000: inst_decode_fn = 9'b0001_xx_xx_0; // BEQ
                        3'b001: inst_decode_fn = 9'b1011_xx_xx_0; // BNE
                        3'b100: inst_decode_fn = 9'b1100_xx_xx_0; // BLT
                        3'b101: inst_decode_fn = 9'b1101_xx_xx_0; // BGE
                        3'b110: inst_decode_fn = 9'b1000_xx_xx_0; // BLTU
                        3'b111: inst_decode_fn = 9'b1001_xx_xx_0; // BGEU
                    
                    endcase
                end
                2'b10: begin // Arithmetic/Logic
                    case (funct3) 
                        3'b000: begin // ADD/SUB
                            if (funct7b5 == 1'b0)
                                inst_decode_fn = 9'b0000_xx_xx_0; // ADD
                            else if (funct7b5 == 1'b1)
                                inst_decode_fn = 9'b0001_xx_xx_0; // SUB
                        end
                        3'b001: inst_decode_fn = 9'b0101_xx_xx_1; // sll
                        3'b010: inst_decode_fn = 9'b1100_xx_xx_0; // SLT signed <
                        3'b011: inst_decode_fn = 9'b1000_xx_xx_0; // SLTU  <
                        3'b100: inst_decode_fn = 9'b0100_xx_xx_0; // XOR
                        3'b101: begin // SRL/SRA
                            if (funct7b5 == 1'b0)
                                inst_decode_fn = 9'b0110_xx_xx_1; // srl
                            else if (funct7b5 == 1'b1)
                                inst_decode_fn = 9'b0111_xx_xx_1; // sra
                        end
                        3'b110: inst_decode_fn = 9'b0011_xx_xx_0; // OR 
                        3'b111: inst_decode_fn = 9'b0010_xx_xx_0; // AND 
                    
                    endcase
                end 
                2'b11: begin // addi (I-type:19系)
                    case (funct3) 
                        3'b000: inst_decode_fn = 9'b0000_xx_xx_x; // ADDI
                        3'b001: inst_decode_fn = 9'b0101_xx_xx_x; // SLLI <<
                        3'b010: inst_decode_fn = 9'b1100_xx_xx_x; // slti : signed <
                        3'b011: inst_decode_fn = 9'b1000_xx_xx_x; // sltiu : <
                        3'b100: inst_decode_fn = 9'b0100_xx_xx_x; // XORI
                        3'b101: begin // SRLI/SRAI
                            if (funct7b5 == 1'b0)
                                inst_decode_fn = 9'b0110_xx_xx_x; // SRLI
                            else if (funct7b5 == 1'b1)
                                inst_decode_fn = 9'b0111_xx_xx_x; // SRAI
                        end
                        3'b110: inst_decode_fn = 9'b0011_xx_xx_x; // ORI
                        3'b111: inst_decode_fn = 9'b0010_xx_xx_x; // ANDI
                    
                    endcase
                end
                default: begin
                    inst_decode_fn = 9'bxxxx_xxxx_x;
                end
            endcase
        end
    endfunction

    assign {alu_ctrl, byte_size, sgn_ext_src, rd2ext_src} = inst_decode_fn(alu_op, funct3, funct7b5);


endmodule

/*    // following code is generated by GPT4.
    always @(alu_op) begin

        // Decode ALU operations
        case (alu_op) 
            2'b00: begin // Load/Store
                case (funct3)
                    3'b000: begin //1byte load/store(lb/sb)
                        alu_ctrl <= 4'b0000; 
                        byte_size <= 2'b10; // this is 1byte l/s
                        sgn_ext_src <= 2'b01; // this is lb
                    end
                    3'b001: begin //2byte load/store(lh/sh)
                        alu_ctrl <= 4'b0000;
                        byte_size <= 2'b01; // this is 2byte l/s
                        sgn_ext_src <= 2'b10; // this is lh
                    end
                    3'b010: begin // ADD (store/load)
                        alu_ctrl <= 4'b0000;
                        byte_size <= 2'b00; // this is 4byte l/s
                    end
                    // lbu(100) , lhu(101)の実装をしていない！
                    // 実装はしたが、lb,lhの符号拡張を自作実装することが発覚したのでその配線追加とモジュール追加。
                    3'b100: begin //1byte load/store(lbu/sbu)
                        alu_ctrl <= 4'b0000; 
                        byte_size <= 2'b10; // this is 1byte l/s
                    end
                    3'b101: begin //2byte load/store(lhu/shu)
                        alu_ctrl <= 4'b0000;
                        byte_size <= 2'b01; // this is 2byte l/s
                    end
                endcase
            end

            2'b01: begin // Branch
                case (funct3)
                    3'b000: alu_ctrl <= 4'b0001; // BEQ (isbranch←1, 引き算後zeroフラグをもらう)
                    3'b001: alu_ctrl <= 4'b1011; // BNE 
                    3'b100: alu_ctrl <= 4'b1100; // BLT 
                    3'b101: alu_ctrl <= 4'b1101; // BGE 
                    3'b110: alu_ctrl <= 4'b1000; // BLTU 
                    3'b111: alu_ctrl <= 4'b1001; // BGEU 
                endcase
            end

            2'b10: begin // Arithmetic/Logic
                case (funct3)
                    3'b000: begin // ADD/SUB
                        if (funct7b5 == 1'b0)
                            alu_ctrl <= 4'b0000; // ADD
                        else if (funct7b5 == 1'b1)
                            alu_ctrl <= 4'b0001; // SUB
                    end

                    3'b001: alu_ctrl <= 4'b0101; // SLL
                    3'b010: alu_ctrl <= 4'b1100; // SLT signed <
                    3'b011: alu_ctrl <= 4'b1000; // SLTU  <
                    3'b100: alu_ctrl <= 4'b0100; // XOR
                    3'b101: begin // SRL/SRA
                        if (funct7b5 == 1'b0)
                            alu_ctrl <= 4'b0110; // srl
                        else if (funct7b5 == 1'b1)
                            alu_ctrl <= 4'b0111; // sra
                    end

                    3'b110: alu_ctrl <= 4'b0011; // OR 
                    3'b111: alu_ctrl <= 4'b0010; // AND 
                endcase
            end
            2'b11: begin // addi (I-type:19系)
                case (funct3)
                    3'b000: alu_ctrl <= 4'b0000; // ADDI
                    3'b001: alu_ctrl <= 4'b0101; // SLLI <<
                    3'b010: alu_ctrl <= 4'b1100; // slti : signed <
                    3'b011: alu_ctrl <= 4'b1000; // sltiu : <
                    3'b100: alu_ctrl <= 4'b0100; // XORI
                    3'b101: begin // SRLI/SRAI
                        if (funct7b5 == 1'b0)
                            alu_ctrl <= 4'b0110; // SRLI
                        else if (funct7b5 == 1'b1)
                            alu_ctrl <= 4'b0111; // SRAI
                    end
                    3'b110: alu_ctrl <= 4'b0011; // ORI
                    3'b111: alu_ctrl <= 4'b0010; // ANDI
                endcase
            end
            default: begin
                alu_ctrl = 4'bxxxx;
            end
        endcase
    end
    */