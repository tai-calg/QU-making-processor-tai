module inst_decoder(
    input [1:0] alu_op,
    input [2:0] funct3,
    input funct7b5,
    output wire [3:0] alu_ctrl,
    output wire [1:0] byte_size,
    output wire [1:0] sgn_ext_src
);


    function [7:0] inst_decode_fn(
        input [1:0] alu_op,
        input [2:0] funct3,
        input funct7b5
    );
        // output = 8'b aluctrl_bytesize_sgnextsrc
        begin
            case (alu_op)
                2'b00: begin // Load
                    case (funct3) 
                        3'b000: inst_decode_fn = 8'b0000_10_01; //1byte load(lb)
                        3'b001: inst_decode_fn = 8'b0000_01_10;//2byte load(lh)
                        3'b010: inst_decode_fn = 8'b0000_00_00; //4byte load(lw)
                        3'b100: inst_decode_fn = 8'b0000_10_00;//1byte load(lbu)
                    endcase
                end
                2'b01: begin // Branch
                    case (funct3) 
                        3'b000: inst_decode_fn = 8'b0001_xx_xx; // BEQ
                        3'b001: inst_decode_fn = 8'b1011_xx_xx; // BNE
                        3'b100: inst_decode_fn = 8'b1100_xx_xx; // BLT
                        3'b101: inst_decode_fn = 8'b1101_xx_xx; // BGE
                        3'b110: inst_decode_fn = 8'b1000_xx_xx; // BLTU
                        3'b111: inst_decode_fn = 8'b1001_xx_xx; // BGEU
                    
                    endcase
                end
                2'b10: begin // Arithmetic/Logic
                    case (funct3) 
                        3'b000: begin // ADD/SUB
                            if (funct7b5 == 1'b0)
                                inst_decode_fn = 8'b0000_xx_xx; // ADD
                            else if (funct7b5 == 1'b1)
                                inst_decode_fn = 8'b0001_xx_xx; // SUB
                        end
                        3'b001: inst_decode_fn = 8'b0101_xx_xx; // SLL
                        3'b010: inst_decode_fn = 8'b1100_xx_xx; // SLT signed <
                        3'b011: inst_decode_fn = 8'b1000_xx_xx; // SLTU  <
                        3'b100: inst_decode_fn = 8'b0100_xx_xx; // XOR
                        3'b101: begin // SRL/SRA
                            if (funct7b5 == 1'b0)
                                inst_decode_fn = 8'b0110_xx_xx; // srl
                            else if (funct7b5 == 1'b1)
                                inst_decode_fn = 8'b0111_xx_xx; // sra
                        end
                        3'b110: inst_decode_fn = 8'b0011_xx_xx; // OR 
                        3'b111: inst_decode_fn = 8'b0010_xx_xx; // AND 
                    
                    endcase
                end 
                2'b11: begin // addi (I-type:19系)
                    case (funct3) 
                        3'b000: inst_decode_fn = 8'b0000_xx_xx; // ADDI
                        3'b001: inst_decode_fn = 8'b0101_xx_xx; // SLLI <<
                        3'b010: inst_decode_fn = 8'b1100_xx_xx; // slti : signed <
                        3'b011: inst_decode_fn = 8'b1000_xx_xx; // sltiu : <
                        3'b100: inst_decode_fn = 8'b0100_xx_xx; // XORI
                        3'b101: begin // SRLI/SRAI
                            if (funct7b5 == 1'b0)
                                inst_decode_fn = 8'b0110_xx_xx; // SRLI
                            else if (funct7b5 == 1'b1)
                                inst_decode_fn = 8'b0111_xx_xx; // SRAI
                        end
                        3'b110: inst_decode_fn = 8'b0011_xx_xx; // ORI
                        3'b111: inst_decode_fn = 8'b0010_xx_xx; // ANDI
                    
                    endcase
                end
                default: begin
                    inst_decode_fn = 8'bxxxx_xxxx;
                end
            endcase
        end
    endfunction

    assign {alu_ctrl, byte_size, sgn_ext_src} = inst_decode_fn(alu_op, funct3, funct7b5);


endmodule

/*    // following code is generated by GPT4.
    always @(alu_op) begin

        // Decode ALU operations
        case (alu_op) 
            2'b00: begin // Load/Store
                case (funct3)
                    3'b000: begin //1byte load/store(lb/sb)
                        alu_ctrl <= 4'b0000; 
                        byte_size <= 2'b10; // this is 1byte l/s
                        sgn_ext_src <= 2'b01; // this is lb
                    end
                    3'b001: begin //2byte load/store(lh/sh)
                        alu_ctrl <= 4'b0000;
                        byte_size <= 2'b01; // this is 2byte l/s
                        sgn_ext_src <= 2'b10; // this is lh
                    end
                    3'b010: begin // ADD (store/load)
                        alu_ctrl <= 4'b0000;
                        byte_size <= 2'b00; // this is 4byte l/s
                    end
                    // lbu(100) , lhu(101)の実装をしていない！
                    //TODO: 実装はしたが、lb,lhの符号拡張を自作実装することが発覚したのでその配線追加とモジュール追加。
                    3'b100: begin //1byte load/store(lbu/sbu)
                        alu_ctrl <= 4'b0000; 
                        byte_size <= 2'b10; // this is 1byte l/s
                    end
                    3'b101: begin //2byte load/store(lhu/shu)
                        alu_ctrl <= 4'b0000;
                        byte_size <= 2'b01; // this is 2byte l/s
                    end
                endcase
            end

            2'b01: begin // Branch
                case (funct3)
                    3'b000: alu_ctrl <= 4'b0001; // BEQ (isbranch←1, 引き算後zeroフラグをもらう)
                    3'b001: alu_ctrl <= 4'b1011; // BNE 
                    3'b100: alu_ctrl <= 4'b1100; // BLT 
                    3'b101: alu_ctrl <= 4'b1101; // BGE 
                    3'b110: alu_ctrl <= 4'b1000; // BLTU 
                    3'b111: alu_ctrl <= 4'b1001; // BGEU 
                endcase
            end

            2'b10: begin // Arithmetic/Logic
                case (funct3)
                    3'b000: begin // ADD/SUB
                        if (funct7b5 == 1'b0)
                            alu_ctrl <= 4'b0000; // ADD
                        else if (funct7b5 == 1'b1)
                            alu_ctrl <= 4'b0001; // SUB
                    end

                    3'b001: alu_ctrl <= 4'b0101; // SLL
                    3'b010: alu_ctrl <= 4'b1100; // SLT signed <
                    3'b011: alu_ctrl <= 4'b1000; // SLTU  <
                    3'b100: alu_ctrl <= 4'b0100; // XOR
                    3'b101: begin // SRL/SRA
                        if (funct7b5 == 1'b0)
                            alu_ctrl <= 4'b0110; // srl
                        else if (funct7b5 == 1'b1)
                            alu_ctrl <= 4'b0111; // sra
                    end

                    3'b110: alu_ctrl <= 4'b0011; // OR 
                    3'b111: alu_ctrl <= 4'b0010; // AND 
                endcase
            end
            2'b11: begin // addi (I-type:19系)
                case (funct3)
                    3'b000: alu_ctrl <= 4'b0000; // ADDI
                    3'b001: alu_ctrl <= 4'b0101; // SLLI <<
                    3'b010: alu_ctrl <= 4'b1100; // slti : signed <
                    3'b011: alu_ctrl <= 4'b1000; // sltiu : <
                    3'b100: alu_ctrl <= 4'b0100; // XORI
                    3'b101: begin // SRLI/SRAI
                        if (funct7b5 == 1'b0)
                            alu_ctrl <= 4'b0110; // SRLI
                        else if (funct7b5 == 1'b1)
                            alu_ctrl <= 4'b0111; // SRAI
                    end
                    3'b110: alu_ctrl <= 4'b0011; // ORI
                    3'b111: alu_ctrl <= 4'b0010; // ANDI
                endcase
            end
            default: begin
                alu_ctrl = 4'bxxxx;
            end
        endcase
    end
    */