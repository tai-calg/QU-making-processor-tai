
module adder(
    input wire [31:0] a,
    input wire [31:0] b,
    output wire [31:0] out,
);
    assign pc_target = pc + immext;
endmodule

